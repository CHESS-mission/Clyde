// ********************************************************************/
// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// SVN Revision Information:
// SVN $Revision: 5996 $
// SVN $Date: 2009-01-16 11:28:16 +0000 (Fri, 16 Jan 2009) $
//
// ********************************************************************/
`timescale 1ns/100ps
module
CoreApbSram_l1I
(
CoreApbSram_lOl
,
CoreApbSram_OIl
,
CoreApbSram_OII
,
CoreApbSram_IIl
,
CoreApbSram_lIl
,
CoreApbSram_Oll
,
CoreApbSram_Ill
,
CoreApbSram_lll
)
;
parameter
CoreApbSram_OOl
=
512
;
localparam
CoreApbSram_O1l
=
1
;
input
[
7
:
0
]
CoreApbSram_lOl
;
input
CoreApbSram_OII
;
input
CoreApbSram_IIl
;
input
[
12
:
0
]
CoreApbSram_lIl
;
input
[
12
:
0
]
CoreApbSram_Oll
;
input
CoreApbSram_Ill
;
input
CoreApbSram_lll
;
output
[
7
:
0
]
CoreApbSram_OIl
;
reg
[
7
:
0
]
CoreApbSram_OIl
;
reg
[
12
:
9
]
CoreApbSram_I1l
;
reg
[
1
:
0
]
CoreApbSram_l1l
;
reg
[
1
:
0
]
CoreApbSram_OO0
;
reg
[
1
:
0
]
CoreApbSram_IO0
;
reg
[
1
:
0
]
CoreApbSram_lO0
;
reg
[
1
:
0
]
CoreApbSram_OI0
;
reg
[
1
:
0
]
CoreApbSram_II0
;
reg
[
1
:
0
]
CoreApbSram_lI0
;
reg
[
1
:
0
]
CoreApbSram_Ol0
;
reg
[
1
:
0
]
CoreApbSram_Il0
;
reg
[
1
:
0
]
CoreApbSram_ll0
;
reg
[
1
:
0
]
CoreApbSram_O00
;
reg
[
1
:
0
]
CoreApbSram_I00
;
reg
[
1
:
0
]
CoreApbSram_l00
;
reg
[
1
:
0
]
CoreApbSram_O10
;
reg
[
1
:
0
]
CoreApbSram_I10
;
reg
[
1
:
0
]
CoreApbSram_l10
;
reg
CoreApbSram_OO1
;
reg
CoreApbSram_IO1
;
reg
CoreApbSram_lO1
;
reg
CoreApbSram_OI1
;
reg
CoreApbSram_II1
;
reg
CoreApbSram_lI1
;
reg
CoreApbSram_Ol1
;
reg
CoreApbSram_Il1
;
reg
CoreApbSram_ll1
;
reg
CoreApbSram_O01
;
reg
CoreApbSram_I01
;
reg
CoreApbSram_l01
;
reg
CoreApbSram_O11
;
reg
CoreApbSram_I11
;
reg
CoreApbSram_l11
;
reg
CoreApbSram_OOOI
;
reg
CoreApbSram_IOOI
;
reg
CoreApbSram_lOOI
;
reg
CoreApbSram_OIOI
;
reg
CoreApbSram_IIOI
;
reg
CoreApbSram_lIOI
;
reg
CoreApbSram_OlOI
;
reg
CoreApbSram_IlOI
;
reg
CoreApbSram_llOI
;
reg
CoreApbSram_O0OI
;
reg
CoreApbSram_I0OI
;
reg
CoreApbSram_l0OI
;
reg
CoreApbSram_O1OI
;
reg
CoreApbSram_I1OI
;
reg
CoreApbSram_l1OI
;
reg
CoreApbSram_OOII
;
reg
CoreApbSram_IOII
;
reg
[
7
:
0
]
CoreApbSram_lOII
;
reg
[
7
:
0
]
CoreApbSram_OIII
;
reg
[
7
:
0
]
CoreApbSram_IIII
;
reg
[
7
:
0
]
CoreApbSram_lIII
;
reg
[
7
:
0
]
CoreApbSram_OlII
;
reg
[
7
:
0
]
CoreApbSram_IlII
;
reg
[
7
:
0
]
CoreApbSram_llII
;
reg
[
7
:
0
]
CoreApbSram_O0II
;
reg
[
7
:
0
]
CoreApbSram_I0II
;
reg
[
7
:
0
]
CoreApbSram_l0II
;
reg
[
7
:
0
]
CoreApbSram_O1II
;
reg
[
7
:
0
]
CoreApbSram_I1II
;
reg
[
7
:
0
]
CoreApbSram_l1II
;
reg
[
7
:
0
]
CoreApbSram_OOlI
;
reg
[
7
:
0
]
CoreApbSram_IOlI
;
reg
[
7
:
0
]
CoreApbSram_lOlI
;
wire
[
7
:
0
]
CoreApbSram_llI
;
wire
[
7
:
0
]
CoreApbSram_IlI
;
wire
[
7
:
0
]
CoreApbSram_OlI
;
wire
[
7
:
0
]
CoreApbSram_lII
;
wire
[
7
:
0
]
CoreApbSram_OIlI
;
wire
[
7
:
0
]
CoreApbSram_IIlI
;
wire
[
7
:
0
]
CoreApbSram_lIlI
;
wire
[
7
:
0
]
CoreApbSram_OllI
;
wire
[
7
:
0
]
CoreApbSram_IllI
;
wire
[
7
:
0
]
CoreApbSram_lllI
;
wire
[
7
:
0
]
CoreApbSram_O0lI
;
wire
[
7
:
0
]
CoreApbSram_I0lI
;
wire
[
7
:
0
]
CoreApbSram_l0lI
;
wire
[
7
:
0
]
CoreApbSram_O1lI
;
wire
[
7
:
0
]
CoreApbSram_I1lI
;
wire
[
7
:
0
]
CoreApbSram_l1lI
;
reg
[
11
:
0
]
CoreApbSram_OO0I
;
reg
[
11
:
0
]
CoreApbSram_IO0I
;
reg
[
11
:
0
]
CoreApbSram_lO0I
;
reg
[
11
:
0
]
CoreApbSram_OI0I
;
reg
[
11
:
0
]
CoreApbSram_II0I
;
reg
[
11
:
0
]
CoreApbSram_lI0I
;
reg
[
11
:
0
]
CoreApbSram_Ol0I
;
reg
[
11
:
0
]
CoreApbSram_Il0I
;
reg
[
11
:
0
]
CoreApbSram_ll0I
;
reg
[
11
:
0
]
CoreApbSram_O00I
;
reg
[
11
:
0
]
CoreApbSram_I00I
;
reg
[
11
:
0
]
CoreApbSram_l00I
;
reg
[
11
:
0
]
CoreApbSram_O10I
;
reg
[
11
:
0
]
CoreApbSram_I10I
;
reg
[
11
:
0
]
CoreApbSram_l10I
;
reg
[
11
:
0
]
CoreApbSram_OO1I
;
reg
[
11
:
0
]
CoreApbSram_IO1I
;
reg
[
11
:
0
]
CoreApbSram_lO1I
;
reg
[
11
:
0
]
CoreApbSram_OI1I
;
reg
[
11
:
0
]
CoreApbSram_II1I
;
reg
[
11
:
0
]
CoreApbSram_lI1I
;
reg
[
11
:
0
]
CoreApbSram_Ol1I
;
reg
[
11
:
0
]
CoreApbSram_Il1I
;
reg
[
11
:
0
]
CoreApbSram_ll1I
;
reg
[
11
:
0
]
CoreApbSram_O01I
;
reg
[
11
:
0
]
CoreApbSram_I01I
;
reg
[
11
:
0
]
CoreApbSram_l01I
;
reg
[
11
:
0
]
CoreApbSram_O11I
;
reg
[
11
:
0
]
CoreApbSram_I11I
;
reg
[
11
:
0
]
CoreApbSram_l11I
;
reg
[
11
:
0
]
CoreApbSram_OOOl
;
reg
[
11
:
0
]
CoreApbSram_IOOl
;
wire
CoreApbSram_O1I
;
wire
CoreApbSram_I1I
;
wire
CoreApbSram_lOOl
;
wire
CoreApbSram_OIOl
;
assign
CoreApbSram_O1I
=
!
CoreApbSram_OII
;
assign
CoreApbSram_I1I
=
!
CoreApbSram_IIl
;
assign
CoreApbSram_lOOl
=
1
'b
1
;
assign
CoreApbSram_OIOl
=
1
'b
0
;
always
@
(
posedge
CoreApbSram_Ill
or
negedge
CoreApbSram_lll
)
begin
if
(
!
CoreApbSram_lll
)
CoreApbSram_I1l
[
12
:
9
]
<=
4
'b
0000
;
else
CoreApbSram_I1l
[
12
:
9
]
<=
CoreApbSram_Oll
[
12
:
9
]
;
end
always
@
(
*
)
begin
CoreApbSram_l1l
=
2
'b
0
;
CoreApbSram_OO0
=
2
'b
0
;
CoreApbSram_IO0
=
2
'b
0
;
CoreApbSram_lO0
=
2
'b
0
;
CoreApbSram_OI0
=
2
'b
0
;
CoreApbSram_II0
=
2
'b
0
;
CoreApbSram_lI0
=
2
'b
0
;
CoreApbSram_Ol0
=
2
'b
0
;
CoreApbSram_Il0
=
2
'b
0
;
CoreApbSram_ll0
=
2
'b
0
;
CoreApbSram_O00
=
2
'b
0
;
CoreApbSram_I00
=
2
'b
0
;
CoreApbSram_l00
=
2
'b
0
;
CoreApbSram_O10
=
2
'b
0
;
CoreApbSram_I10
=
2
'b
0
;
CoreApbSram_l10
=
2
'b
0
;
CoreApbSram_OO1
=
1
'b
1
;
CoreApbSram_IO1
=
1
'b
1
;
CoreApbSram_lO1
=
1
'b
1
;
CoreApbSram_OI1
=
1
'b
1
;
CoreApbSram_II1
=
1
'b
1
;
CoreApbSram_lI1
=
1
'b
1
;
CoreApbSram_Ol1
=
1
'b
1
;
CoreApbSram_Il1
=
1
'b
1
;
CoreApbSram_ll1
=
1
'b
1
;
CoreApbSram_O01
=
1
'b
1
;
CoreApbSram_I01
=
1
'b
1
;
CoreApbSram_l01
=
1
'b
1
;
CoreApbSram_O11
=
1
'b
1
;
CoreApbSram_I11
=
1
'b
1
;
CoreApbSram_l11
=
1
'b
1
;
CoreApbSram_OOOI
=
1
'b
1
;
CoreApbSram_IOOI
=
1
'b
1
;
CoreApbSram_lOOI
=
1
'b
1
;
CoreApbSram_OIOI
=
1
'b
1
;
CoreApbSram_IIOI
=
1
'b
1
;
CoreApbSram_lIOI
=
1
'b
1
;
CoreApbSram_OlOI
=
1
'b
1
;
CoreApbSram_IlOI
=
1
'b
1
;
CoreApbSram_llOI
=
1
'b
1
;
CoreApbSram_O0OI
=
1
'b
1
;
CoreApbSram_I0OI
=
1
'b
1
;
CoreApbSram_l0OI
=
1
'b
1
;
CoreApbSram_O1OI
=
1
'b
1
;
CoreApbSram_I1OI
=
1
'b
1
;
CoreApbSram_l1OI
=
1
'b
1
;
CoreApbSram_OOII
=
1
'b
1
;
CoreApbSram_IOII
=
1
'b
1
;
CoreApbSram_lOII
=
8
'b
0
;
CoreApbSram_OIII
=
8
'b
0
;
CoreApbSram_IIII
=
8
'b
0
;
CoreApbSram_lIII
=
8
'b
0
;
CoreApbSram_OlII
=
8
'b
0
;
CoreApbSram_IlII
=
8
'b
0
;
CoreApbSram_llII
=
8
'b
0
;
CoreApbSram_O0II
=
8
'b
0
;
CoreApbSram_I0II
=
8
'b
0
;
CoreApbSram_l0II
=
8
'b
0
;
CoreApbSram_O1II
=
8
'b
0
;
CoreApbSram_I1II
=
8
'b
0
;
CoreApbSram_l1II
=
8
'b
0
;
CoreApbSram_OOlI
=
8
'b
0
;
CoreApbSram_IOlI
=
8
'b
0
;
CoreApbSram_lOlI
=
8
'b
0
;
CoreApbSram_OO0I
=
12
'b
0
;
CoreApbSram_IO0I
=
12
'b
0
;
CoreApbSram_lO0I
=
12
'b
0
;
CoreApbSram_OI0I
=
12
'b
0
;
CoreApbSram_II0I
=
12
'b
0
;
CoreApbSram_lI0I
=
12
'b
0
;
CoreApbSram_Ol0I
=
12
'b
0
;
CoreApbSram_Il0I
=
12
'b
0
;
CoreApbSram_ll0I
=
12
'b
0
;
CoreApbSram_O00I
=
12
'b
0
;
CoreApbSram_I00I
=
12
'b
0
;
CoreApbSram_l00I
=
12
'b
0
;
CoreApbSram_O10I
=
12
'b
0
;
CoreApbSram_I10I
=
12
'b
0
;
CoreApbSram_l10I
=
12
'b
0
;
CoreApbSram_OO1I
=
12
'b
0
;
CoreApbSram_IO1I
=
12
'b
0
;
CoreApbSram_lO1I
=
12
'b
0
;
CoreApbSram_OI1I
=
12
'b
0
;
CoreApbSram_II1I
=
12
'b
0
;
CoreApbSram_lI1I
=
12
'b
0
;
CoreApbSram_Ol1I
=
12
'b
0
;
CoreApbSram_Il1I
=
12
'b
0
;
CoreApbSram_ll1I
=
12
'b
0
;
CoreApbSram_O01I
=
12
'b
0
;
CoreApbSram_I01I
=
12
'b
0
;
CoreApbSram_l01I
=
12
'b
0
;
CoreApbSram_O11I
=
12
'b
0
;
CoreApbSram_I11I
=
12
'b
0
;
CoreApbSram_l11I
=
12
'b
0
;
CoreApbSram_OOOl
=
12
'b
0
;
CoreApbSram_IOOl
=
12
'b
0
;
case
(
CoreApbSram_OOl
)
512
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OO1
=
CoreApbSram_O1I
;
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
CoreApbSram_OIl
=
CoreApbSram_llI
;
end
1024
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
9
]
)
1
'b
0
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
1
'b
1
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
9
]
)
1
'b
0
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
1
'b
1
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
9
]
)
1
'b
0
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
1
'b
1
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
end
endcase
1536
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
2
'b
01
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
2
'b
10
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
2
'b
11
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
2
'b
01
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
2
'b
10
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
2
'b
11
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
2
'b
01
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
2
'b
10
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
2
'b
11
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
10
:
9
]
)
2
'b
00
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
2
'b
01
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
2
'b
10
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
2
'b
11
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
10
:
9
]
)
2
'b
00
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
2
'b
01
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
2
'b
10
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
2
'b
11
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
2
'b
01
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
2
'b
10
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
2
'b
11
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
endcase
end
endcase
2048
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
2
'b
01
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
2
'b
10
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
2
'b
11
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
2
'b
01
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
2
'b
10
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
2
'b
11
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
2
'b
01
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
2
'b
10
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
2
'b
11
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
10
:
9
]
)
2
'b
00
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
2
'b
01
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
2
'b
10
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
2
'b
11
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
10
:
9
]
)
2
'b
00
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
2
'b
01
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
2
'b
10
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
2
'b
11
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
10
:
9
]
)
2
'b
00
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
2
'b
01
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
2
'b
10
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
2
'b
11
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
end
endcase
2560
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
3
'b
001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
3
'b
010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
3
'b
110
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
111
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
3
'b
001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
3
'b
010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
3
'b
110
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
111
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
3
'b
001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
3
'b
010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
111
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
endcase
end
endcase
3072
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
3
'b
001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
3
'b
010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
3
'b
110
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
111
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
3
'b
001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
3
'b
010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
3
'b
110
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
111
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
3
'b
001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
3
'b
010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
111
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
endcase
end
endcase
3584
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
3
'b
001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
3
'b
010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
3
'b
110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
3
'b
111
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
3
'b
001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
3
'b
010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
3
'b
110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
3
'b
111
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
3
'b
001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
3
'b
010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
3
'b
111
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
3
'b
111
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
3
'b
111
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
endcase
end
endcase
4096
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
3
'b
001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
3
'b
010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
3
'b
011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
3
'b
100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
3
'b
101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
3
'b
110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
3
'b
111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
3
'b
001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
3
'b
010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
3
'b
011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
3
'b
100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
3
'b
101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
3
'b
110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
3
'b
111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
3
'b
001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
3
'b
010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
3
'b
011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
3
'b
100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
3
'b
101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
3
'b
110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
3
'b
111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
case
(
CoreApbSram_lIl
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
3
'b
111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
11
:
9
]
)
3
'b
000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
3
'b
111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
11
:
9
]
)
3
'b
000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
3
'b
111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
4608
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
5120
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
5632
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
6144
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_I00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
CoreApbSram_I1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_l01
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_O1OI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_I0lI
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
10
;
CoreApbSram_I00
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_I1II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
6656
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_I00
=
2
'b
11
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
CoreApbSram_I1II
=
CoreApbSram_lOl
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_l01
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_O1OI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_I0lI
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
10
;
CoreApbSram_I00
=
2
'b
10
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_I1II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
7168
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_I00
=
2
'b
11
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_O10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
CoreApbSram_I1II
=
CoreApbSram_lOl
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
CoreApbSram_OOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_l01
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_I11
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_O1OI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_l1OI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_I0lI
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_O1lI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
10
;
CoreApbSram_I00
=
2
'b
10
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_I1II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
7680
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_I00
=
2
'b
11
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_O10
=
2
'b
11
;
CoreApbSram_I10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
CoreApbSram_I1II
=
CoreApbSram_lOl
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
CoreApbSram_OOlI
=
CoreApbSram_lOl
;
CoreApbSram_IOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_l01
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_I11
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_l11
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_O1OI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_l1OI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_OOII
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_I0lI
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_O1lI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_I1lI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
10
;
CoreApbSram_I00
=
2
'b
10
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_I10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_I1II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
CoreApbSram_l11
=
CoreApbSram_O1I
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
CoreApbSram_OOII
=
CoreApbSram_I1I
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_I1lI
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_I10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
CoreApbSram_l11
=
CoreApbSram_O1I
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
CoreApbSram_OOII
=
CoreApbSram_I1I
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_I1lI
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_I10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
CoreApbSram_l11
=
CoreApbSram_O1I
;
4
'b
1111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
CoreApbSram_OOII
=
CoreApbSram_I1I
;
4
'b
1111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_I1lI
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
endcase
end
endcase
default
:
case
(
CoreApbSram_O1l
)
8
:
begin
CoreApbSram_l1l
=
2
'b
11
;
CoreApbSram_OO0
=
2
'b
11
;
CoreApbSram_IO0
=
2
'b
11
;
CoreApbSram_lO0
=
2
'b
11
;
CoreApbSram_OI0
=
2
'b
11
;
CoreApbSram_II0
=
2
'b
11
;
CoreApbSram_lI0
=
2
'b
11
;
CoreApbSram_Ol0
=
2
'b
11
;
CoreApbSram_Il0
=
2
'b
11
;
CoreApbSram_ll0
=
2
'b
11
;
CoreApbSram_O00
=
2
'b
11
;
CoreApbSram_I00
=
2
'b
11
;
CoreApbSram_l00
=
2
'b
11
;
CoreApbSram_O10
=
2
'b
11
;
CoreApbSram_I10
=
2
'b
11
;
CoreApbSram_l10
=
2
'b
11
;
CoreApbSram_OO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lO0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_II0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_lI0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Ol0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_Il0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_ll0I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l00I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_O10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_I10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_l10I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_OO1I
=
{
3
'b
0
,
CoreApbSram_lIl
[
8
:
0
]
}
;
CoreApbSram_IO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lO1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_II1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lI1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Ol1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_Il1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_ll1I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l01I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_O11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_I11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_l11I
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_OOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_IOOl
=
{
3
'b
0
,
CoreApbSram_Oll
[
8
:
0
]
}
;
CoreApbSram_lOII
=
CoreApbSram_lOl
;
CoreApbSram_OIII
=
CoreApbSram_lOl
;
CoreApbSram_IIII
=
CoreApbSram_lOl
;
CoreApbSram_lIII
=
CoreApbSram_lOl
;
CoreApbSram_OlII
=
CoreApbSram_lOl
;
CoreApbSram_IlII
=
CoreApbSram_lOl
;
CoreApbSram_llII
=
CoreApbSram_lOl
;
CoreApbSram_O0II
=
CoreApbSram_lOl
;
CoreApbSram_I0II
=
CoreApbSram_lOl
;
CoreApbSram_l0II
=
CoreApbSram_lOl
;
CoreApbSram_O1II
=
CoreApbSram_lOl
;
CoreApbSram_I1II
=
CoreApbSram_lOl
;
CoreApbSram_l1II
=
CoreApbSram_lOl
;
CoreApbSram_OOlI
=
CoreApbSram_lOl
;
CoreApbSram_IOlI
=
CoreApbSram_lOl
;
CoreApbSram_lOlI
=
CoreApbSram_lOl
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OO1
=
CoreApbSram_O1I
;
4
'b
0001
:
CoreApbSram_IO1
=
CoreApbSram_O1I
;
4
'b
0010
:
CoreApbSram_lO1
=
CoreApbSram_O1I
;
4
'b
0011
:
CoreApbSram_OI1
=
CoreApbSram_O1I
;
4
'b
0100
:
CoreApbSram_II1
=
CoreApbSram_O1I
;
4
'b
0101
:
CoreApbSram_lI1
=
CoreApbSram_O1I
;
4
'b
0110
:
CoreApbSram_Ol1
=
CoreApbSram_O1I
;
4
'b
0111
:
CoreApbSram_Il1
=
CoreApbSram_O1I
;
4
'b
1000
:
CoreApbSram_ll1
=
CoreApbSram_O1I
;
4
'b
1001
:
CoreApbSram_O01
=
CoreApbSram_O1I
;
4
'b
1010
:
CoreApbSram_I01
=
CoreApbSram_O1I
;
4
'b
1011
:
CoreApbSram_l01
=
CoreApbSram_O1I
;
4
'b
1100
:
CoreApbSram_O11
=
CoreApbSram_O1I
;
4
'b
1101
:
CoreApbSram_I11
=
CoreApbSram_O1I
;
4
'b
1110
:
CoreApbSram_l11
=
CoreApbSram_O1I
;
4
'b
1111
:
CoreApbSram_OOOI
=
CoreApbSram_O1I
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_IOOI
=
CoreApbSram_I1I
;
4
'b
0001
:
CoreApbSram_lOOI
=
CoreApbSram_I1I
;
4
'b
0010
:
CoreApbSram_OIOI
=
CoreApbSram_I1I
;
4
'b
0011
:
CoreApbSram_IIOI
=
CoreApbSram_I1I
;
4
'b
0100
:
CoreApbSram_lIOI
=
CoreApbSram_I1I
;
4
'b
0101
:
CoreApbSram_OlOI
=
CoreApbSram_I1I
;
4
'b
0110
:
CoreApbSram_IlOI
=
CoreApbSram_I1I
;
4
'b
0111
:
CoreApbSram_llOI
=
CoreApbSram_I1I
;
4
'b
1000
:
CoreApbSram_O0OI
=
CoreApbSram_I1I
;
4
'b
1001
:
CoreApbSram_I0OI
=
CoreApbSram_I1I
;
4
'b
1010
:
CoreApbSram_l0OI
=
CoreApbSram_I1I
;
4
'b
1011
:
CoreApbSram_O1OI
=
CoreApbSram_I1I
;
4
'b
1100
:
CoreApbSram_I1OI
=
CoreApbSram_I1I
;
4
'b
1101
:
CoreApbSram_l1OI
=
CoreApbSram_I1I
;
4
'b
1110
:
CoreApbSram_OOII
=
CoreApbSram_I1I
;
4
'b
1111
:
CoreApbSram_IOII
=
CoreApbSram_I1I
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
CoreApbSram_llI
;
4
'b
0001
:
CoreApbSram_OIl
=
CoreApbSram_IlI
;
4
'b
0010
:
CoreApbSram_OIl
=
CoreApbSram_OlI
;
4
'b
0011
:
CoreApbSram_OIl
=
CoreApbSram_lII
;
4
'b
0100
:
CoreApbSram_OIl
=
CoreApbSram_OIlI
;
4
'b
0101
:
CoreApbSram_OIl
=
CoreApbSram_IIlI
;
4
'b
0110
:
CoreApbSram_OIl
=
CoreApbSram_lIlI
;
4
'b
0111
:
CoreApbSram_OIl
=
CoreApbSram_OllI
;
4
'b
1000
:
CoreApbSram_OIl
=
CoreApbSram_IllI
;
4
'b
1001
:
CoreApbSram_OIl
=
CoreApbSram_lllI
;
4
'b
1010
:
CoreApbSram_OIl
=
CoreApbSram_O0lI
;
4
'b
1011
:
CoreApbSram_OIl
=
CoreApbSram_I0lI
;
4
'b
1100
:
CoreApbSram_OIl
=
CoreApbSram_l0lI
;
4
'b
1101
:
CoreApbSram_OIl
=
CoreApbSram_O1lI
;
4
'b
1110
:
CoreApbSram_OIl
=
CoreApbSram_I1lI
;
4
'b
1111
:
CoreApbSram_OIl
=
CoreApbSram_l1lI
;
endcase
end
4
:
begin
CoreApbSram_l1l
=
2
'b
10
;
CoreApbSram_OO0
=
2
'b
10
;
CoreApbSram_IO0
=
2
'b
10
;
CoreApbSram_lO0
=
2
'b
10
;
CoreApbSram_OI0
=
2
'b
10
;
CoreApbSram_II0
=
2
'b
10
;
CoreApbSram_lI0
=
2
'b
10
;
CoreApbSram_Ol0
=
2
'b
10
;
CoreApbSram_Il0
=
2
'b
10
;
CoreApbSram_ll0
=
2
'b
10
;
CoreApbSram_O00
=
2
'b
10
;
CoreApbSram_I00
=
2
'b
10
;
CoreApbSram_l00
=
2
'b
10
;
CoreApbSram_O10
=
2
'b
10
;
CoreApbSram_I10
=
2
'b
10
;
CoreApbSram_l10
=
2
'b
10
;
CoreApbSram_OO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lO0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_II0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_lI0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Ol0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_Il0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_ll0I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l00I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_O10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_I10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_l10I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_OO1I
=
{
2
'b
0
,
CoreApbSram_lIl
[
9
:
0
]
}
;
CoreApbSram_IO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lO1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_II1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lI1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Ol1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_Il1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_ll1I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l01I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_O11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_I11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_l11I
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_OOOl
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_IOOl
=
{
2
'b
0
,
CoreApbSram_Oll
[
9
:
0
]
}
;
CoreApbSram_lOII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IIII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lIII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_OlII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_IlII
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_llII
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_O0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_I0II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_l0II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_O1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_I1II
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_l1II
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_OOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
CoreApbSram_IOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
3
:
0
]
;
CoreApbSram_lOlI
[
3
:
0
]
=
CoreApbSram_lOl
[
7
:
4
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_IlI
[
3
:
0
]
,
CoreApbSram_llI
[
3
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
3
:
0
]
,
CoreApbSram_OlI
[
3
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_IIlI
[
3
:
0
]
,
CoreApbSram_OIlI
[
3
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
3
:
0
]
,
CoreApbSram_lIlI
[
3
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_lllI
[
3
:
0
]
,
CoreApbSram_IllI
[
3
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
3
:
0
]
,
CoreApbSram_O0lI
[
3
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_O1lI
[
3
:
0
]
,
CoreApbSram_l0lI
[
3
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
3
:
0
]
,
CoreApbSram_I1lI
[
3
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
3
:
0
]
,
CoreApbSram_I1lI
[
3
:
0
]
}
;
endcase
end
2
:
begin
CoreApbSram_l1l
=
2
'b
01
;
CoreApbSram_OO0
=
2
'b
01
;
CoreApbSram_IO0
=
2
'b
01
;
CoreApbSram_lO0
=
2
'b
01
;
CoreApbSram_OI0
=
2
'b
01
;
CoreApbSram_II0
=
2
'b
01
;
CoreApbSram_lI0
=
2
'b
01
;
CoreApbSram_Ol0
=
2
'b
01
;
CoreApbSram_Il0
=
2
'b
01
;
CoreApbSram_ll0
=
2
'b
01
;
CoreApbSram_O00
=
2
'b
01
;
CoreApbSram_I00
=
2
'b
01
;
CoreApbSram_l00
=
2
'b
01
;
CoreApbSram_O10
=
2
'b
01
;
CoreApbSram_I10
=
2
'b
01
;
CoreApbSram_l10
=
2
'b
01
;
CoreApbSram_OO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lO0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_II0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_lI0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Ol0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_Il0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_ll0I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l00I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_O10I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_I10I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_l10I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_OO1I
=
{
1
'b
0
,
CoreApbSram_lIl
[
10
:
0
]
}
;
CoreApbSram_IO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lO1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_II1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lI1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Ol1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_Il1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_ll1I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l01I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_O11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_I11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_l11I
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_OOOl
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_IOOl
=
{
1
'b
0
,
CoreApbSram_Oll
[
10
:
0
]
}
;
CoreApbSram_lOII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OIII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IIII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lIII
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_OlII
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_IlII
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_llII
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_O0II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_I0II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_l0II
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_O1II
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_I1II
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
CoreApbSram_l1II
[
1
:
0
]
=
CoreApbSram_lOl
[
1
:
0
]
;
CoreApbSram_OOlI
[
1
:
0
]
=
CoreApbSram_lOl
[
3
:
2
]
;
CoreApbSram_IOlI
[
1
:
0
]
=
CoreApbSram_lOl
[
5
:
4
]
;
CoreApbSram_lOlI
[
1
:
0
]
=
CoreApbSram_lOl
[
7
:
6
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_lII
[
1
:
0
]
,
CoreApbSram_OlI
[
1
:
0
]
,
CoreApbSram_IlI
[
1
:
0
]
,
CoreApbSram_llI
[
1
:
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
1
:
0
]
,
CoreApbSram_lIlI
[
1
:
0
]
,
CoreApbSram_IIlI
[
1
:
0
]
,
CoreApbSram_OIlI
[
1
:
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_I0lI
[
1
:
0
]
,
CoreApbSram_O0lI
[
1
:
0
]
,
CoreApbSram_lllI
[
1
:
0
]
,
CoreApbSram_IllI
[
1
:
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
1
:
0
]
,
CoreApbSram_I1lI
[
1
:
0
]
,
CoreApbSram_O1lI
[
1
:
0
]
,
CoreApbSram_l0lI
[
1
:
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
1
:
0
]
,
CoreApbSram_I1lI
[
1
:
0
]
,
CoreApbSram_O1lI
[
1
:
0
]
,
CoreApbSram_l0lI
[
1
:
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
1
:
0
]
,
CoreApbSram_I1lI
[
1
:
0
]
,
CoreApbSram_O1lI
[
1
:
0
]
,
CoreApbSram_l0lI
[
1
:
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
1
:
0
]
,
CoreApbSram_I1lI
[
1
:
0
]
,
CoreApbSram_O1lI
[
1
:
0
]
,
CoreApbSram_l0lI
[
1
:
0
]
}
;
endcase
end
default
:
begin
CoreApbSram_l1l
=
2
'b
00
;
CoreApbSram_OO0
=
2
'b
00
;
CoreApbSram_IO0
=
2
'b
00
;
CoreApbSram_lO0
=
2
'b
00
;
CoreApbSram_OI0
=
2
'b
00
;
CoreApbSram_II0
=
2
'b
00
;
CoreApbSram_lI0
=
2
'b
00
;
CoreApbSram_Ol0
=
2
'b
00
;
CoreApbSram_Il0
=
2
'b
00
;
CoreApbSram_ll0
=
2
'b
00
;
CoreApbSram_O00
=
2
'b
00
;
CoreApbSram_I00
=
2
'b
00
;
CoreApbSram_l00
=
2
'b
00
;
CoreApbSram_O10
=
2
'b
00
;
CoreApbSram_I10
=
2
'b
00
;
CoreApbSram_l10
=
2
'b
00
;
CoreApbSram_OO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lO0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_II0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_lI0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Ol0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_Il0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_ll0I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_O00I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_I00I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_l00I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_O10I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_I10I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_l10I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_OO1I
=
{
CoreApbSram_lIl
[
11
:
0
]
}
;
CoreApbSram_IO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lO1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_II1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lI1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Ol1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_Il1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_ll1I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O01I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_I01I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_l01I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_O11I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_I11I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_l11I
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_OOOl
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_IOOl
=
{
CoreApbSram_Oll
[
11
:
0
]
}
;
CoreApbSram_lOII
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_OIII
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_IIII
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_lIII
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_OlII
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_IlII
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_llII
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_O0II
[
0
]
=
CoreApbSram_lOl
[
7
]
;
CoreApbSram_I0II
[
0
]
=
CoreApbSram_lOl
[
0
]
;
CoreApbSram_l0II
[
0
]
=
CoreApbSram_lOl
[
1
]
;
CoreApbSram_O1II
[
0
]
=
CoreApbSram_lOl
[
2
]
;
CoreApbSram_I1II
[
0
]
=
CoreApbSram_lOl
[
3
]
;
CoreApbSram_l1II
[
0
]
=
CoreApbSram_lOl
[
4
]
;
CoreApbSram_OOlI
[
0
]
=
CoreApbSram_lOl
[
5
]
;
CoreApbSram_IOlI
[
0
]
=
CoreApbSram_lOl
[
6
]
;
CoreApbSram_lOlI
[
0
]
=
CoreApbSram_lOl
[
7
]
;
case
(
CoreApbSram_lIl
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0001
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0010
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0011
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0100
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0101
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0110
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
0111
:
{
CoreApbSram_Il1
,
CoreApbSram_Ol1
,
CoreApbSram_lI1
,
CoreApbSram_II1
,
CoreApbSram_OI1
,
CoreApbSram_lO1
,
CoreApbSram_IO1
,
CoreApbSram_OO1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1000
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1001
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1010
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1011
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1100
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1101
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1110
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
4
'b
1111
:
{
CoreApbSram_OOOI
,
CoreApbSram_l11
,
CoreApbSram_I11
,
CoreApbSram_O11
,
CoreApbSram_l01
,
CoreApbSram_I01
,
CoreApbSram_O01
,
CoreApbSram_ll1
}
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
endcase
case
(
CoreApbSram_Oll
[
12
:
9
]
)
4
'b
0000
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0001
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0010
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0011
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0100
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0101
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0110
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
0111
:
{
CoreApbSram_llOI
,
CoreApbSram_IlOI
,
CoreApbSram_OlOI
,
CoreApbSram_lIOI
,
CoreApbSram_IIOI
,
CoreApbSram_OIOI
,
CoreApbSram_lOOI
,
CoreApbSram_IOOI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1000
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1001
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1010
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1011
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1100
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1101
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1110
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
4
'b
1111
:
{
CoreApbSram_IOII
,
CoreApbSram_OOII
,
CoreApbSram_l1OI
,
CoreApbSram_I1OI
,
CoreApbSram_O1OI
,
CoreApbSram_l0OI
,
CoreApbSram_I0OI
,
CoreApbSram_O0OI
}
=
{
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
,
CoreApbSram_I1I
}
;
endcase
case
(
CoreApbSram_I1l
[
12
:
9
]
)
4
'b
0000
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0001
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0010
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0011
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0100
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0101
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0110
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
0111
:
CoreApbSram_OIl
=
{
CoreApbSram_OllI
[
0
]
,
CoreApbSram_lIlI
[
0
]
,
CoreApbSram_IIlI
[
0
]
,
CoreApbSram_OIlI
[
0
]
,
CoreApbSram_lII
[
0
]
,
CoreApbSram_OlI
[
0
]
,
CoreApbSram_IlI
[
0
]
,
CoreApbSram_llI
[
0
]
}
;
4
'b
1000
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1001
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1010
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1011
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1100
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1101
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1110
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
4
'b
1111
:
CoreApbSram_OIl
=
{
CoreApbSram_l1lI
[
0
]
,
CoreApbSram_I1lI
[
0
]
,
CoreApbSram_O1lI
[
0
]
,
CoreApbSram_l0lI
[
0
]
,
CoreApbSram_I0lI
[
0
]
,
CoreApbSram_O0lI
[
0
]
,
CoreApbSram_lllI
[
0
]
,
CoreApbSram_IllI
[
0
]
}
;
endcase
end
endcase
endcase
end
RAM4K9
CoreApbSram_IIOl
(
.ADDRA11
(
CoreApbSram_OO0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_IO1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_OO0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_IO1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_OO0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_IO1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_OO0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_IO1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_OO0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_IO1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_OO0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_IO1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_OO0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_IO1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_OO0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_IO1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_OO0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_IO1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_OO0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_IO1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_OO0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_IO1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_OO0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_IO1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_lOII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_lOII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_lOII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_lOII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_lOII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_lOII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_lOII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_lOII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_llI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_llI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_llI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_llI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_llI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_llI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_llI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_llI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_l1l
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_l1l
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_l1l
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_l1l
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_OO1
)
,
.BLKB
(
CoreApbSram_IOOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_lIOl
(
.ADDRA11
(
CoreApbSram_IO0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_lO1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_IO0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_lO1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_IO0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_lO1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_IO0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_lO1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_IO0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_lO1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_IO0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_lO1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_IO0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_lO1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_IO0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_lO1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_IO0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_lO1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_IO0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_lO1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_IO0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_lO1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_IO0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_lO1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_OIII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_OIII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_OIII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_OIII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_OIII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_OIII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_OIII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_OIII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_IlI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_IlI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_IlI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_IlI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_IlI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_IlI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_IlI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_IlI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_OO0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_OO0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_OO0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_OO0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_IO1
)
,
.BLKB
(
CoreApbSram_lOOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_OlOl
(
.ADDRA11
(
CoreApbSram_lO0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_OI1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_lO0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_OI1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_lO0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_OI1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_lO0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_OI1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_lO0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_OI1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_lO0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_OI1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_lO0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_OI1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_lO0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_OI1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_lO0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_OI1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_lO0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_OI1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_lO0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_OI1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_lO0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_OI1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_IIII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_IIII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_IIII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_IIII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_IIII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_IIII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_IIII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_IIII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_OlI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_OlI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_OlI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_OlI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_OlI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_OlI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_OlI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_OlI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_IO0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_IO0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_IO0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_IO0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_lO1
)
,
.BLKB
(
CoreApbSram_OIOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_IlOl
(
.ADDRA11
(
CoreApbSram_OI0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_II1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_OI0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_II1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_OI0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_II1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_OI0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_II1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_OI0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_II1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_OI0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_II1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_OI0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_II1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_OI0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_II1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_OI0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_II1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_OI0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_II1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_OI0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_II1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_OI0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_II1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_lIII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_lIII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_lIII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_lIII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_lIII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_lIII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_lIII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_lIII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_lII
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_lII
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_lII
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_lII
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_lII
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_lII
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_lII
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_lII
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_lO0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_lO0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_lO0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_lO0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_OI1
)
,
.BLKB
(
CoreApbSram_IIOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_llOl
(
.ADDRA11
(
CoreApbSram_II0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_lI1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_II0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_lI1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_II0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_lI1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_II0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_lI1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_II0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_lI1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_II0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_lI1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_II0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_lI1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_II0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_lI1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_II0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_lI1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_II0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_lI1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_II0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_lI1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_II0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_lI1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_OlII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_OlII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_OlII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_OlII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_OlII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_OlII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_OlII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_OlII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_OIlI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_OIlI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_OIlI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_OIlI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_OIlI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_OIlI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_OIlI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_OIlI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_OI0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_OI0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_OI0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_OI0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_II1
)
,
.BLKB
(
CoreApbSram_lIOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_O0Ol
(
.ADDRA11
(
CoreApbSram_lI0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_Ol1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_lI0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_Ol1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_lI0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_Ol1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_lI0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_Ol1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_lI0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_Ol1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_lI0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_Ol1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_lI0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_Ol1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_lI0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_Ol1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_lI0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_Ol1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_lI0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_Ol1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_lI0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_Ol1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_lI0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_Ol1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_IlII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_IlII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_IlII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_IlII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_IlII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_IlII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_IlII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_IlII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_IIlI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_IIlI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_IIlI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_IIlI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_IIlI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_IIlI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_IIlI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_IIlI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_II0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_II0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_II0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_II0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_lI1
)
,
.BLKB
(
CoreApbSram_OlOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_I0Ol
(
.ADDRA11
(
CoreApbSram_Ol0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_Il1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_Ol0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_Il1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_Ol0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_Il1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_Ol0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_Il1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_Ol0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_Il1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_Ol0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_Il1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_Ol0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_Il1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_Ol0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_Il1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_Ol0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_Il1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_Ol0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_Il1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_Ol0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_Il1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_Ol0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_Il1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_llII
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_llII
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_llII
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_llII
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_llII
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_llII
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_llII
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_llII
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_lIlI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_lIlI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_lIlI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_lIlI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_lIlI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_lIlI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_lIlI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_lIlI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_lI0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_lI0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_lI0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_lI0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_Ol1
)
,
.BLKB
(
CoreApbSram_IlOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_l0Ol
(
.ADDRA11
(
CoreApbSram_Il0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_ll1I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_Il0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_ll1I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_Il0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_ll1I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_Il0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_ll1I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_Il0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_ll1I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_Il0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_ll1I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_Il0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_ll1I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_Il0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_ll1I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_Il0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_ll1I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_Il0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_ll1I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_Il0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_ll1I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_Il0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_ll1I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_O0II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_O0II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_O0II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_O0II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_O0II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_O0II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_O0II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_O0II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_OllI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_OllI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_OllI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_OllI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_OllI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_OllI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_OllI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_OllI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_Ol0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_Ol0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_Ol0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_Ol0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_Il1
)
,
.BLKB
(
CoreApbSram_llOI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_O1Ol
(
.ADDRA11
(
CoreApbSram_ll0I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_O01I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_ll0I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_O01I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_ll0I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_O01I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_ll0I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_O01I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_ll0I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_O01I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_ll0I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_O01I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_ll0I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_O01I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_ll0I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_O01I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_ll0I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_O01I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_ll0I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_O01I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_ll0I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_O01I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_ll0I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_O01I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_I0II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_I0II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_I0II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_I0II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_I0II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_I0II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_I0II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_I0II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_IllI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_IllI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_IllI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_IllI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_IllI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_IllI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_IllI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_IllI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_Il0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_Il0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_Il0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_Il0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_ll1
)
,
.BLKB
(
CoreApbSram_O0OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_I1Ol
(
.ADDRA11
(
CoreApbSram_O00I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_I01I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_O00I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_I01I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_O00I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_I01I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_O00I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_I01I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_O00I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_I01I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_O00I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_I01I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_O00I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_I01I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_O00I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_I01I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_O00I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_I01I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_O00I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_I01I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_O00I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_I01I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_O00I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_I01I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_l0II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_l0II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_l0II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_l0II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_l0II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_l0II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_l0II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_l0II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_lllI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_lllI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_lllI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_lllI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_lllI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_lllI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_lllI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_lllI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_ll0
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_ll0
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_ll0
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_ll0
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_O01
)
,
.BLKB
(
CoreApbSram_I0OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_l1Ol
(
.ADDRA11
(
CoreApbSram_I00I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_l01I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_I00I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_l01I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_I00I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_l01I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_I00I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_l01I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_I00I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_l01I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_I00I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_l01I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_I00I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_l01I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_I00I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_l01I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_I00I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_l01I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_I00I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_l01I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_I00I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_l01I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_I00I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_l01I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_O1II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_O1II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_O1II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_O1II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_O1II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_O1II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_O1II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_O1II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_O0lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_O0lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_O0lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_O0lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_O0lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_O0lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_O0lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_O0lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_O00
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_O00
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_O00
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_O00
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_I01
)
,
.BLKB
(
CoreApbSram_l0OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_OOIl
(
.ADDRA11
(
CoreApbSram_l00I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_O11I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_l00I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_O11I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_l00I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_O11I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_l00I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_O11I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_l00I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_O11I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_l00I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_O11I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_l00I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_O11I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_l00I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_O11I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_l00I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_O11I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_l00I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_O11I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_l00I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_O11I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_l00I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_O11I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_I1II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_I1II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_I1II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_I1II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_I1II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_I1II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_I1II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_I1II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_I0lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_I0lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_I0lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_I0lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_I0lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_I0lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_I0lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_I0lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_I00
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_I00
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_I00
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_I00
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_l01
)
,
.BLKB
(
CoreApbSram_O1OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_IOIl
(
.ADDRA11
(
CoreApbSram_O10I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_I11I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_O10I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_I11I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_O10I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_I11I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_O10I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_I11I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_O10I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_I11I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_O10I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_I11I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_O10I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_I11I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_O10I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_I11I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_O10I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_I11I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_O10I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_I11I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_O10I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_I11I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_O10I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_I11I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_l1II
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_l1II
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_l1II
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_l1II
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_l1II
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_l1II
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_l1II
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_l1II
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_l0lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_l0lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_l0lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_l0lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_l0lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_l0lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_l0lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_l0lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_l00
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_l00
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_l00
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_l00
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_O11
)
,
.BLKB
(
CoreApbSram_I1OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_lOIl
(
.ADDRA11
(
CoreApbSram_I10I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_l11I
[
11
]
)
,
.ADDRA10
(
CoreApbSram_I10I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_l11I
[
10
]
)
,
.ADDRA9
(
CoreApbSram_I10I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_l11I
[
9
]
)
,
.ADDRA8
(
CoreApbSram_I10I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_l11I
[
8
]
)
,
.ADDRA7
(
CoreApbSram_I10I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_l11I
[
7
]
)
,
.ADDRA6
(
CoreApbSram_I10I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_l11I
[
6
]
)
,
.ADDRA5
(
CoreApbSram_I10I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_l11I
[
5
]
)
,
.ADDRA4
(
CoreApbSram_I10I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_l11I
[
4
]
)
,
.ADDRA3
(
CoreApbSram_I10I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_l11I
[
3
]
)
,
.ADDRA2
(
CoreApbSram_I10I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_l11I
[
2
]
)
,
.ADDRA1
(
CoreApbSram_I10I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_l11I
[
1
]
)
,
.ADDRA0
(
CoreApbSram_I10I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_l11I
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_OOlI
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_OOlI
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_OOlI
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_OOlI
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_OOlI
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_OOlI
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_OOlI
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_OOlI
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_O1lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_O1lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_O1lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_O1lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_O1lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_O1lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_O1lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_O1lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_O10
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_O10
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_O10
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_O10
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_I11
)
,
.BLKB
(
CoreApbSram_l1OI
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_OIIl
(
.ADDRA11
(
CoreApbSram_l10I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_OOOl
[
11
]
)
,
.ADDRA10
(
CoreApbSram_l10I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_OOOl
[
10
]
)
,
.ADDRA9
(
CoreApbSram_l10I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_OOOl
[
9
]
)
,
.ADDRA8
(
CoreApbSram_l10I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_OOOl
[
8
]
)
,
.ADDRA7
(
CoreApbSram_l10I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_OOOl
[
7
]
)
,
.ADDRA6
(
CoreApbSram_l10I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_OOOl
[
6
]
)
,
.ADDRA5
(
CoreApbSram_l10I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_OOOl
[
5
]
)
,
.ADDRA4
(
CoreApbSram_l10I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_OOOl
[
4
]
)
,
.ADDRA3
(
CoreApbSram_l10I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_OOOl
[
3
]
)
,
.ADDRA2
(
CoreApbSram_l10I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_OOOl
[
2
]
)
,
.ADDRA1
(
CoreApbSram_l10I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_OOOl
[
1
]
)
,
.ADDRA0
(
CoreApbSram_l10I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_OOOl
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_IOlI
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_IOlI
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_IOlI
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_IOlI
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_IOlI
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_IOlI
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_IOlI
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_IOlI
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_I1lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_I1lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_I1lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_I1lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_I1lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_I1lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_I1lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_I1lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_I10
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_I10
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_I10
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_I10
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_l11
)
,
.BLKB
(
CoreApbSram_OOII
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
RAM4K9
CoreApbSram_IIIl
(
.ADDRA11
(
CoreApbSram_OO1I
[
11
]
)
,
.ADDRB11
(
CoreApbSram_IOOl
[
11
]
)
,
.ADDRA10
(
CoreApbSram_OO1I
[
10
]
)
,
.ADDRB10
(
CoreApbSram_IOOl
[
10
]
)
,
.ADDRA9
(
CoreApbSram_OO1I
[
9
]
)
,
.ADDRB9
(
CoreApbSram_IOOl
[
9
]
)
,
.ADDRA8
(
CoreApbSram_OO1I
[
8
]
)
,
.ADDRB8
(
CoreApbSram_IOOl
[
8
]
)
,
.ADDRA7
(
CoreApbSram_OO1I
[
7
]
)
,
.ADDRB7
(
CoreApbSram_IOOl
[
7
]
)
,
.ADDRA6
(
CoreApbSram_OO1I
[
6
]
)
,
.ADDRB6
(
CoreApbSram_IOOl
[
6
]
)
,
.ADDRA5
(
CoreApbSram_OO1I
[
5
]
)
,
.ADDRB5
(
CoreApbSram_IOOl
[
5
]
)
,
.ADDRA4
(
CoreApbSram_OO1I
[
4
]
)
,
.ADDRB4
(
CoreApbSram_IOOl
[
4
]
)
,
.ADDRA3
(
CoreApbSram_OO1I
[
3
]
)
,
.ADDRB3
(
CoreApbSram_IOOl
[
3
]
)
,
.ADDRA2
(
CoreApbSram_OO1I
[
2
]
)
,
.ADDRB2
(
CoreApbSram_IOOl
[
2
]
)
,
.ADDRA1
(
CoreApbSram_OO1I
[
1
]
)
,
.ADDRB1
(
CoreApbSram_IOOl
[
1
]
)
,
.ADDRA0
(
CoreApbSram_OO1I
[
0
]
)
,
.ADDRB0
(
CoreApbSram_IOOl
[
0
]
)
,
.DINA8
(
CoreApbSram_OIOl
)
,
.DINB8
(
CoreApbSram_OIOl
)
,
.DINA7
(
CoreApbSram_lOlI
[
7
]
)
,
.DINB7
(
CoreApbSram_OIOl
)
,
.DINA6
(
CoreApbSram_lOlI
[
6
]
)
,
.DINB6
(
CoreApbSram_OIOl
)
,
.DINA5
(
CoreApbSram_lOlI
[
5
]
)
,
.DINB5
(
CoreApbSram_OIOl
)
,
.DINA4
(
CoreApbSram_lOlI
[
4
]
)
,
.DINB4
(
CoreApbSram_OIOl
)
,
.DINA3
(
CoreApbSram_lOlI
[
3
]
)
,
.DINB3
(
CoreApbSram_OIOl
)
,
.DINA2
(
CoreApbSram_lOlI
[
2
]
)
,
.DINB2
(
CoreApbSram_OIOl
)
,
.DINA1
(
CoreApbSram_lOlI
[
1
]
)
,
.DINB1
(
CoreApbSram_OIOl
)
,
.DINA0
(
CoreApbSram_lOlI
[
0
]
)
,
.DINB0
(
CoreApbSram_OIOl
)
,
.DOUTA8
(
)
,
.DOUTB8
(
)
,
.DOUTA7
(
)
,
.DOUTB7
(
CoreApbSram_l1lI
[
7
]
)
,
.DOUTA6
(
)
,
.DOUTB6
(
CoreApbSram_l1lI
[
6
]
)
,
.DOUTA5
(
)
,
.DOUTB5
(
CoreApbSram_l1lI
[
5
]
)
,
.DOUTA4
(
)
,
.DOUTB4
(
CoreApbSram_l1lI
[
4
]
)
,
.DOUTA3
(
)
,
.DOUTB3
(
CoreApbSram_l1lI
[
3
]
)
,
.DOUTA2
(
)
,
.DOUTB2
(
CoreApbSram_l1lI
[
2
]
)
,
.DOUTA1
(
)
,
.DOUTB1
(
CoreApbSram_l1lI
[
1
]
)
,
.DOUTA0
(
)
,
.DOUTB0
(
CoreApbSram_l1lI
[
0
]
)
,
.WIDTHA1
(
CoreApbSram_l10
[
1
]
)
,
.WIDTHB1
(
CoreApbSram_l10
[
1
]
)
,
.WIDTHA0
(
CoreApbSram_l10
[
0
]
)
,
.WIDTHB0
(
CoreApbSram_l10
[
0
]
)
,
.PIPEA
(
CoreApbSram_OIOl
)
,
.PIPEB
(
CoreApbSram_OIOl
)
,
.WMODEA
(
CoreApbSram_OIOl
)
,
.WMODEB
(
CoreApbSram_OIOl
)
,
.BLKA
(
CoreApbSram_OOOI
)
,
.BLKB
(
CoreApbSram_IOII
)
,
.WENA
(
CoreApbSram_OIOl
)
,
.WENB
(
CoreApbSram_lOOl
)
,
.CLKA
(
CoreApbSram_Ill
)
,
.CLKB
(
CoreApbSram_Ill
)
,
.RESET
(
CoreApbSram_lll
)
)
;
endmodule
