// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/100ps
module
Minimal_SoC_CoreUARTapb_0_fifo_256x8
(
CUARTOOOI
,
CUARTIOOI
,
CUARTlOOI
,
CUARTOIOI
,
WRB
,
RDB
,
RESET
,
FULL
,
EMPTY
)
;
output
[
7
:
0
]
CUARTOOOI
;
input
CUARTIOOI
;
input
CUARTlOOI
;
input
[
7
:
0
]
CUARTOIOI
;
input
WRB
;
input
RDB
;
input
RESET
;
output
FULL
;
output
EMPTY
;
parameter
SYNC_RESET
=
0
;
parameter
[
7
:
0
]
CUARTOIlI
=
255
;
wire
AEMPTY
,
AFULL
,
FULL
,
EMPTY
;
reg
[
7
:
0
]
CUARTOOOI
;
wire
[
7
:
0
]
CUARTl00I
;
always
@
(
posedge
CUARTIOOI
)
begin
CUARTOOOI
<=
CUARTl00I
;
end
Minimal_SoC_CoreUARTapb_0_fifo_256x8_pa3
Minimal_SoC_CoreUARTapb_0_fifo_256x8_pa3
(
.CUARTIIOl
(
CUARTOIOI
)
,
.CUARTlI1I
(
CUARTl00I
)
,
.CUARTll1I
(
WRB
)
,
.CUARTO01I
(
RDB
)
,
.CUARTlOOI
(
CUARTlOOI
)
,
.CUARTIOOI
(
CUARTIOOI
)
,
.AEMPTY
(
AEMPTY
)
,
.AFULL
(
GEQTH
)
,
.FULL
(
FULL
)
,
.EMPTY
(
EMPTY
)
,
.RESET
(
RESET
)
,
.CUARTOIlI
(
CUARTOIlI
)
)
;
endmodule
module
Minimal_SoC_CoreUARTapb_0_fifo_256x8_pa3
(
CUARTIIOl
,
CUARTlI1I
,
CUARTll1I
,
CUARTO01I
,
CUARTlOOI
,
CUARTIOOI
,
FULL
,
EMPTY
,
RESET
,
AEMPTY
,
AFULL
,
CUARTOIlI
)
;
input
[
7
:
0
]
CUARTIIOl
;
output
[
7
:
0
]
CUARTlI1I
;
input
CUARTll1I
,
CUARTO01I
,
CUARTlOOI
,
CUARTIOOI
;
output
FULL
,
EMPTY
;
input
RESET
;
output
AEMPTY
,
AFULL
;
input
[
7
:
0
]
CUARTOIlI
;
wire
CUARTlIOl
,
VCC
,
GND
;
VCC
CUARTl11I
(
.Y
(
VCC
)
)
;
GND
CUARTOOOl
(
.Y
(
GND
)
)
;
INV
CUARTOlOl
(
.A
(
CUARTO01I
)
,
.Y
(
CUARTlIOl
)
)
;
FIFO4K18
CUARTIlOl
(
.AEVAL11
(
GND
)
,
.AEVAL10
(
GND
)
,
.AEVAL9
(
GND
)
,
.AEVAL8
(
GND
)
,
.AEVAL7
(
GND
)
,
.AEVAL6
(
GND
)
,
.AEVAL5
(
GND
)
,
.AEVAL4
(
GND
)
,
.AEVAL3
(
VCC
)
,
.AEVAL2
(
GND
)
,
.AEVAL1
(
GND
)
,
.AEVAL0
(
GND
)
,
.AFVAL11
(
GND
)
,
.AFVAL10
(
CUARTOIlI
[
7
]
)
,
.AFVAL9
(
CUARTOIlI
[
6
]
)
,
.AFVAL8
(
CUARTOIlI
[
5
]
)
,
.AFVAL7
(
CUARTOIlI
[
4
]
)
,
.AFVAL6
(
CUARTOIlI
[
3
]
)
,
.AFVAL5
(
CUARTOIlI
[
2
]
)
,
.AFVAL4
(
CUARTOIlI
[
1
]
)
,
.AFVAL3
(
CUARTOIlI
[
0
]
)
,
.AFVAL2
(
GND
)
,
.AFVAL1
(
GND
)
,
.AFVAL0
(
GND
)
,
.WD17
(
GND
)
,
.WD16
(
GND
)
,
.WD15
(
GND
)
,
.WD14
(
GND
)
,
.WD13
(
GND
)
,
.WD12
(
GND
)
,
.WD11
(
GND
)
,
.WD10
(
GND
)
,
.WD9
(
GND
)
,
.WD8
(
GND
)
,
.WD7
(
CUARTIIOl
[
7
]
)
,
.WD6
(
CUARTIIOl
[
6
]
)
,
.WD5
(
CUARTIIOl
[
5
]
)
,
.WD4
(
CUARTIIOl
[
4
]
)
,
.WD3
(
CUARTIIOl
[
3
]
)
,
.WD2
(
CUARTIIOl
[
2
]
)
,
.WD1
(
CUARTIIOl
[
1
]
)
,
.WD0
(
CUARTIIOl
[
0
]
)
,
.WW0
(
VCC
)
,
.WW1
(
VCC
)
,
.WW2
(
GND
)
,
.RW0
(
VCC
)
,
.RW1
(
VCC
)
,
.RW2
(
GND
)
,
.RPIPE
(
GND
)
,
.WEN
(
CUARTll1I
)
,
.REN
(
CUARTlIOl
)
,
.WBLK
(
GND
)
,
.RBLK
(
GND
)
,
.WCLK
(
CUARTlOOI
)
,
.RCLK
(
CUARTIOOI
)
,
.RESET
(
RESET
)
,
.ESTOP
(
VCC
)
,
.FSTOP
(
VCC
)
,
.RD17
(
)
,
.RD16
(
)
,
.RD15
(
)
,
.RD14
(
)
,
.RD13
(
)
,
.RD12
(
)
,
.RD11
(
)
,
.RD10
(
)
,
.RD9
(
)
,
.RD8
(
)
,
.RD7
(
CUARTlI1I
[
7
]
)
,
.RD6
(
CUARTlI1I
[
6
]
)
,
.RD5
(
CUARTlI1I
[
5
]
)
,
.RD4
(
CUARTlI1I
[
4
]
)
,
.RD3
(
CUARTlI1I
[
3
]
)
,
.RD2
(
CUARTlI1I
[
2
]
)
,
.RD1
(
CUARTlI1I
[
1
]
)
,
.RD0
(
CUARTlI1I
[
0
]
)
,
.FULL
(
)
,
.AFULL
(
FULL
)
,
.EMPTY
(
EMPTY
)
,
.AEMPTY
(
AEMPTY
)
)
;
endmodule
