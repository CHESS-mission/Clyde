// ********************************************************************/
// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// SVN Revision Information:
// SVN $Revision: 5996 $
// SVN $Date: 2009-01-16 11:28:16 +0000 (Fri, 16 Jan 2009) $
//
// ********************************************************************/
`timescale 1ns/100ps
module
COREAPBSRAM
(
	PCLK
,
PRESETN
,
	PSEL
,
PENABLE
,
PWRITE
,
PADDR
,
PWDATA
,
PRDATA
,
PSLVERR
,
PREADY
)
;
parameter
FAMILY
=
17
;
parameter
APB_DWIDTH
=
32
;
parameter
NUM_LOCATIONS_DWIDTH32
=
512
;
parameter
NUM_LOCATIONS_DWIDTH24
=
512
;
parameter
NUM_LOCATIONS_DWIDTH16
=
512
;
parameter
NUM_LOCATIONS_DWIDTH08
=
512
;
parameter
ADDR_SCHEME
=
0
;
localparam
CoreApbSram_O
=
NUM_LOCATIONS_DWIDTH32
;
localparam
CoreApbSram_I
=
NUM_LOCATIONS_DWIDTH24
;
localparam
CoreApbSram_l
=
CoreApbSram_OI
(
NUM_LOCATIONS_DWIDTH16
)
;
localparam
CoreApbSram_II
=
CoreApbSram_lI
(
NUM_LOCATIONS_DWIDTH16
)
;
localparam
CoreApbSram_Ol
=
CoreApbSram_Il
(
NUM_LOCATIONS_DWIDTH08
)
;
localparam
CoreApbSram_ll
=
CoreApbSram_O0
(
NUM_LOCATIONS_DWIDTH08
)
;
localparam
CoreApbSram_I0
=
CoreApbSram_l0
(
NUM_LOCATIONS_DWIDTH08
)
;
localparam
CoreApbSram_O1
=
CoreApbSram_I1
(
NUM_LOCATIONS_DWIDTH08
)
;
localparam
CoreApbSram_l1
=
(
CoreApbSram_II
==
0
)
?
512
:
CoreApbSram_II
;
localparam
CoreApbSram_OOI
=
(
CoreApbSram_ll
==
0
)
?
512
:
CoreApbSram_ll
;
localparam
CoreApbSram_IOI
=
(
CoreApbSram_I0
==
0
)
?
512
:
CoreApbSram_I0
;
localparam
CoreApbSram_lOI
=
(
CoreApbSram_O1
==
0
)
?
512
:
CoreApbSram_O1
;
input
	PCLK
;
input
PRESETN
;
input
	PSEL
;
input
PENABLE
;
input
PWRITE
;
input
[
16
:
0
]
PADDR
;
input
[
APB_DWIDTH
-
1
:
0
]
PWDATA
;
output
reg
[
APB_DWIDTH
-
1
:
0
]
PRDATA
;
output
PSLVERR
;
output
PREADY
;
reg
[
3
:
0
]
CoreApbSram_OII
;
reg
[
12
:
0
]
CoreApbSram_III
;
wire
[
7
:
0
]
CoreApbSram_lII
;
wire
[
7
:
0
]
CoreApbSram_OlI
;
wire
[
7
:
0
]
CoreApbSram_IlI
;
wire
[
7
:
0
]
CoreApbSram_llI
;
wire
[
7
:
0
]
CoreApbSram_O0I
;
wire
[
7
:
0
]
CoreApbSram_I0I
;
wire
[
7
:
0
]
CoreApbSram_l0I
;
wire
CoreApbSram_O1I
;
wire
CoreApbSram_I1I
;
function
[
31
:
0
]
CoreApbSram_OI
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH16
;
begin
if
(
NUM_LOCATIONS_DWIDTH16
<
8193
)
begin
CoreApbSram_OI
=
NUM_LOCATIONS_DWIDTH16
;
end
else
begin
CoreApbSram_OI
=
8192
;
end
end
endfunction
function
[
31
:
0
]
CoreApbSram_lI
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH16
;
begin
if
(
NUM_LOCATIONS_DWIDTH16
<
8193
)
begin
CoreApbSram_lI
=
0
;
end
else
begin
CoreApbSram_lI
=
NUM_LOCATIONS_DWIDTH16
-
8192
;
end
end
endfunction
function
[
31
:
0
]
CoreApbSram_Il
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH08
;
begin
if
(
NUM_LOCATIONS_DWIDTH08
<
8193
)
begin
CoreApbSram_Il
=
NUM_LOCATIONS_DWIDTH08
;
end
else
begin
CoreApbSram_Il
=
8192
;
end
end
endfunction
function
[
31
:
0
]
CoreApbSram_O0
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH08
;
begin
if
(
NUM_LOCATIONS_DWIDTH08
<
8193
)
begin
CoreApbSram_O0
=
0
;
end
else
if
(
NUM_LOCATIONS_DWIDTH08
>
8192
&&
NUM_LOCATIONS_DWIDTH08
<
16385
)
begin
CoreApbSram_O0
=
NUM_LOCATIONS_DWIDTH08
-
8192
;
end
else
begin
CoreApbSram_O0
=
8192
;
end
end
endfunction
function
[
31
:
0
]
CoreApbSram_l0
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH08
;
begin
if
(
NUM_LOCATIONS_DWIDTH08
<
16385
)
begin
CoreApbSram_l0
=
0
;
end
else
if
(
NUM_LOCATIONS_DWIDTH08
>
16384
&&
NUM_LOCATIONS_DWIDTH08
<
24577
)
begin
CoreApbSram_l0
=
NUM_LOCATIONS_DWIDTH08
-
16384
;
end
else
begin
CoreApbSram_l0
=
8192
;
end
end
endfunction
function
[
31
:
0
]
CoreApbSram_I1
;
input
[
31
:
0
]
NUM_LOCATIONS_DWIDTH08
;
begin
if
(
NUM_LOCATIONS_DWIDTH08
<
24577
)
begin
CoreApbSram_I1
=
0
;
end
else
begin
CoreApbSram_I1
=
NUM_LOCATIONS_DWIDTH08
-
24576
;
end
end
endfunction
assign
PSLVERR
=
1
'b
0
;
assign
PREADY
=
1
'b
1
;
assign
CoreApbSram_O1I
=
PWRITE
&&
PENABLE
&&
	PSEL
;
assign
CoreApbSram_I1I
=
~
PWRITE
&&
~
PENABLE
&&
	PSEL
;
generate
if
(
APB_DWIDTH
==
32
)
begin
always
@
(
*
)
begin
case
(
ADDR_SCHEME
)
1
:
begin
CoreApbSram_III
=
PADDR
[
12
:
0
]
;
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_lII
,
CoreApbSram_OlI
,
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
end
default
:
begin
CoreApbSram_III
=
PADDR
[
14
:
2
]
;
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_lII
,
CoreApbSram_OlI
,
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
end
endcase
end
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_O
)
)
CoreApbSram_IOl
(
.CoreApbSram_lOl
(
PWDATA
[
31
:
24
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_lII
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
3
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_O
)
)
CoreApbSram_O0l
(
.CoreApbSram_lOl
(
PWDATA
[
23
:
16
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_OlI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
2
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_O
)
)
CoreApbSram_I0l
(
.CoreApbSram_lOl
(
PWDATA
[
15
:
8
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_IlI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
1
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_O
)
)
CoreApbSram_l0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_llI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
0
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
end
else
if
(
APB_DWIDTH
==
24
)
begin
always
@
(
*
)
begin
case
(
ADDR_SCHEME
)
1
:
begin
CoreApbSram_III
=
PADDR
[
12
:
0
]
;
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_OlI
,
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
end
default
:
begin
CoreApbSram_III
=
PADDR
[
14
:
2
]
;
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
CoreApbSram_O1I
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_OlI
,
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
end
endcase
end
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_I
)
)
CoreApbSram_O0l
(
.CoreApbSram_lOl
(
PWDATA
[
23
:
16
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_OlI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
2
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_I
)
)
CoreApbSram_I0l
(
.CoreApbSram_lOl
(
PWDATA
[
15
:
8
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_IlI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
1
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_I
)
)
CoreApbSram_l0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_llI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
0
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
end
else
if
(
APB_DWIDTH
==
16
)
begin
always
@
(
*
)
begin
case
(
ADDR_SCHEME
)
1
:
begin
CoreApbSram_III
=
PADDR
[
12
:
0
]
;
case
(
PADDR
[
13
]
)
1
'b
0
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
1
'b
1
:
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
}
;
default
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
endcase
case
(
PADDR
[
13
]
)
1
'b
0
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
1
'b
1
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_lII
,
CoreApbSram_OlI
}
;
default
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
endcase
end
default
:
begin
CoreApbSram_III
=
PADDR
[
14
:
2
]
;
case
(
PADDR
[
15
]
)
1
'b
0
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
,
CoreApbSram_O1I
}
;
1
'b
1
:
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
}
;
default
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
endcase
case
(
PADDR
[
15
]
)
1
'b
0
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
1
'b
1
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_lII
,
CoreApbSram_OlI
}
;
default
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
{
CoreApbSram_IlI
,
CoreApbSram_llI
}
;
endcase
end
endcase
end
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_l1
)
)
CoreApbSram_IOl
(
.CoreApbSram_lOl
(
PWDATA
[
15
:
8
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_O0I
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
3
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_l1
)
)
CoreApbSram_O0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_I0I
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
2
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_l
)
)
CoreApbSram_I0l
(
.CoreApbSram_lOl
(
PWDATA
[
15
:
8
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_IlI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
1
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_l
)
)
CoreApbSram_l0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_llI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
0
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
assign
CoreApbSram_lII
=
(
CoreApbSram_II
==
0
)
?
8
'b
0
:
CoreApbSram_O0I
;
assign
CoreApbSram_OlI
=
(
CoreApbSram_II
==
0
)
?
8
'b
0
:
CoreApbSram_I0I
;
end
else
begin
always
@
(
*
)
begin
case
(
ADDR_SCHEME
)
1
:
begin
CoreApbSram_III
=
PADDR
[
12
:
0
]
;
case
(
PADDR
[
14
:
13
]
)
2
'b
00
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
}
;
2
'b
01
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
,
1
'b
0
}
;
2
'b
10
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
}
;
2
'b
11
:
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
default
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
endcase
case
(
PADDR
[
14
:
13
]
)
2
'b
00
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_llI
;
2
'b
01
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_IlI
;
2
'b
10
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_OlI
;
2
'b
11
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_lII
;
default
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_llI
;
endcase
end
default
:
begin
CoreApbSram_III
=
PADDR
[
14
:
2
]
;
case
(
PADDR
[
16
:
15
]
)
2
'b
00
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
}
;
2
'b
01
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
CoreApbSram_O1I
,
1
'b
0
}
;
2
'b
10
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
}
;
2
'b
11
:
CoreApbSram_OII
[
3
:
0
]
=
{
CoreApbSram_O1I
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
default
:
CoreApbSram_OII
[
3
:
0
]
=
{
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
;
endcase
case
(
PADDR
[
16
:
15
]
)
2
'b
00
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_llI
;
2
'b
01
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_IlI
;
2
'b
10
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_OlI
;
2
'b
11
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_lII
;
default
:
PRDATA
[
APB_DWIDTH
-
1
:
0
]
=
CoreApbSram_llI
;
endcase
end
endcase
end
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_lOI
)
)
CoreApbSram_IOl
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_O0I
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
3
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_IOI
)
)
CoreApbSram_O0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_I0I
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
2
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_OOI
)
)
CoreApbSram_I0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_l0I
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
1
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
CoreApbSram_l1I
#
(
.CoreApbSram_OOl
(
CoreApbSram_Ol
)
)
CoreApbSram_l0l
(
.CoreApbSram_lOl
(
PWDATA
[
7
:
0
]
)
,
.CoreApbSram_OIl
(
CoreApbSram_llI
)
,
.CoreApbSram_OII
(
CoreApbSram_OII
[
0
]
)
,
.CoreApbSram_IIl
(
CoreApbSram_I1I
)
,
.CoreApbSram_lIl
(
CoreApbSram_III
)
,
.CoreApbSram_Oll
(
CoreApbSram_III
)
,
.CoreApbSram_Ill
(
	PCLK
)
,
.CoreApbSram_lll
(
PRESETN
)
)
;
assign
CoreApbSram_lII
=
(
CoreApbSram_O1
==
0
)
?
8
'b
0
:
CoreApbSram_O0I
;
assign
CoreApbSram_OlI
=
(
CoreApbSram_I0
==
0
)
?
8
'b
0
:
CoreApbSram_I0I
;
assign
CoreApbSram_IlI
=
(
CoreApbSram_ll
==
0
)
?
8
'b
0
:
CoreApbSram_l0I
;
end
endgenerate
endmodule
